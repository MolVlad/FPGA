module top(
    input CLK,
    input TXD,
	 input S2,
	 
	 output RXD,
    output DS_EN1, DS_EN2, DS_EN3, DS_EN4,
    output DS_A, DS_B, DS_C, DS_D, DS_E, DS_F, DS_G, DS_DP
);

/* -------------- Clock ------------------ */

wire uart_clk;

custome_clk_div #(.x(18), .y(1250)) custome_clk_div(.clk(CLK), .clk_out(uart_clk));	// 1250 * 38400 = 48.000.000

/* -------------- UART TX ---------------- */

wire [7:0]uart_data;
wire flag_complete;

uart_in uart_in(.clk(uart_clk), .in(TXD), .data(uart_data), .flag_complete(flag_complete));

/* -------------- Display ---------------- */

wire [15:0]data;

wire [3:0]hex_data;

ascii_to_hex ascii_to_hex(.ascii(uart_data), .hex(hex_data));

display_shift display_shift(.clk(flag_complete), .num(hex_data), .data(data));

wire [3:0]anodes;
assign {DS_EN1, DS_EN2, DS_EN3, DS_EN4} = ~anodes;

wire [7:0]seg;
assign {DS_A, DS_B, DS_C, DS_D, DS_E, DS_F, DS_G, DS_DP} = seg;

hex_display hex_display(.clk(CLK), .data(data), .anodes(anodes), .seg(seg));

/* -------------- UART RX ---------------- */

wire [7:0]ascii;

hex_to_ascii hex_to_ascii(.hex(data[3:0]), .ascii(ascii));

wire uart_in_edge;

posedge_impulse posedge_impulse(.clk(uart_clk), .in(flag_complete), .out(uart_in_edge));

uart_out uart_out(.clk(uart_clk), .data(ascii), .out(RXD), .flag_start(uart_in_edge));

endmodule
